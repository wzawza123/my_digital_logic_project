module pc1 
(
    input i_CLK,
    input i_RST,
    output reg o_CLK
);
    
endmodule