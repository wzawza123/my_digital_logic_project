module pc2
(
    input i_CLK,
    input i_RST,
    output reg o_CLK
);
    initial begin
        o_CLK = 0;
    end

endmodule